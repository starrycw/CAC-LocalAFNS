//
//  1.MODULES:
//
//  1.1 adder_fxx: 
//      ���������xxλ쳲�������ϵ�ļӷ�����
//      ��adder_f05��λǡ�ÿ��Լ���f3+f4=f5
//      Adder_fxx(FNS_n-2_in, FNS_n-1_in, FNS_n_out, FNS_n-1_out, f_flag)
//  
//  1.2 FNSadders_x_y:
//      FNS Adders������en_flag�ļ����·������xΪ����TSV����yΪ����TSV����    
//
//  1.3 coder_x_y, dec_x_y:
//      ���������FTF��������xΪ����TSV����yΪ����TSV����
//
//  1.4 CACcoder_x, CACdec_x:
//      FNS-CAC���������FTF��������xΪλ����
//
// 
//  2.SIMULATION:
//
//  2.1 Simu_x_y:
//      ������֤������xΪ����TSV��Ŀ��yΪ����TSV��Ŀ��
//      ��֤���ݰ�������1���������������ֵ�Ƿ�����������������ֵ����2�������Ƿ�����������������Ѿ�������λ���⣬����λ������FTF������
//      test01:�޹��������
//      test02:����1��ʧЧTSV
//      test03:����2��ʧЧTSV
//      test04:���ڶ��ʧЧTSV������1�������Ϊ������Ŀ��
//      
//  2.2 Simu_x:
//        FNS-CAC�Ĺ�����֤������xΪ����TSV��Ŀ��
//        Ϊ�˼������Ƿ��д���
//        ��֤����1���������������ֵ�Ƿ�����������������ֵ����2�������Ƿ����FTF����